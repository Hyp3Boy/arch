`timescale 1ns / 1ps

module mux8_tb();

reg a0,a1,a2,a3,a4,a5,a6,a7,s0,s1,s2;
wire y;

mux8 m0(a0,a1,a2,a3,a4,a5,a6,a7,s0,s1,s2,y);

initial begin
  $dumpfile("mux8_tb.vcd");
  $dumpvars(0,mux8_tb);
  $monitor("a0=%b a1=%b a2=%b a3=%b a4=%b a5=%b a6=%b a7=%b s0=%b s1=%b s2=%b y=%b",a0,a1,a2,a3,a4,a5,a6,a7,s0,s1,s2,y);
  a0 = 0; a1 = 0; a2 = 0; a3 = 0; a4 = 0; a5 = 0; a6 = 0; a7 = 0; s0 = 0; s1 = 0; s2 = 0;
  #10 a0=0; a1=0; a2=0; a3=0; a4=0; a5=0; a6=0; a7=0; s0=0; s1=0; s2=0;
  #10 a0=0; a1=0; a2=0; a3=0; a4=0; a5=0; a6=0; a7=0; s0=0; s1=0; s2=1;
  #10 a0=0; a1=0; a2=0; a3=0; a4=0; a5=0; a6=0; a7=0; s0=0; s1=1; s2=0;
  #10 a0=0; a1=0; a2=0; a3=0; a4=0; a5=0; a6=0; a7=0; s0=0; s1=1; s2=1;
  #10 a0=0; a1=0; a2=0; a3=0; a4=0; a5=0; a6=0; a7=0; s0=1; s1=0; s2=0;
  #10 a0=0; a1=0; a2=0; a3=0; a4=0; a5=0; a6=0; a7=0; s0=1; s1=0; s2=1;
  #10 a0=0; a1=0; a2=0; a3=0; a4=0; a5=0; a6=0; a7=0; s0=1; s1=1; s2=0;
  #10 a0=0; a1=0; a2=0; a3=0; a4=0; a5=0; a6=0; a7=0; s0=1; s1=1; s2=1;
  #10 a0=0; a1=0; a2=0; a3=0; a4=0; a5=0; a6=0; a7=1; s0=0; s1=0; s2=0;
  #10 a0=0; a1=0; a2=0; a3=0; a4=0; a5=0; a6=0; a7=1; s0=0; s1=0; s2=1;
  #10 a0=0; a1=0; a2=0; a3=0; a4=0; a5=0; a6=0; a7=1; s0=0; s1=1; s2=0;
  #10 a0=0; a1=0; a2=0; a3=0; a4=0; a5=0; a6=0; a7=1; s0=0; s1=1; s2=1;
  #10 a0=0; a1=0; a2=0; a3=0; a4=0; a5=0; a6=0; a7=1; s0=1; s1=0; s2=0;
  #10 a0=0; a1=0; a2=0; a3=0; a4=0; a5=0; a6=0; a7=1; s0=1; s1=0; s2=1;
  #10 a0=0; a1=0; a2=0; a3=0; a4=0; a5=0; a6=0; a7=1; s0=1; s1=1; s2=0;
  #10 a0=0; a1=0; a2=0; a3=0; a4=0; a5=0; a6
=0; a7=1; s0=1; s1=1; s2=1;
  #10 $finish;

end

endmodule

